isa18_2021_2022@localhost.localdomain.32016:1630289278