wackoz@wT14.419742:1640081599