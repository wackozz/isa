isa18_2021_2022@localhost.localdomain.17787:1630289278